module Instruction_memory(
                        
endmodule
